module Lab4_1(F, A);
input [0:3] A;
output [0:1] F;
reg [0:1] F;

always @ (A)
	case(A)
	4'b0000: F[0:1]=2'b00;
	4'b0001: F[0:1]=2'b10;
	4'b0010: F[0:1]=2'b01;
	4'b0011: F[0:1]=2'b11;
	4'b0100: F[0:1]=2'b01;
	4'b0101: F[0:1]=2'b00;
	4'b0110: F[0:1]=2'b10;
	4'b0111: F[0:1]=2'b10;
	4'b1000: F <= 2'b10;
	4'b1001: F <= 2'b10;
	4'b1010: F <= 2'b11;
	4'b1011: F <= 2'b11;
	4'b1100: F <= 2'b11;
	4'b1101: F <= 2'b10;
	4'b1110: F <= 2'b10;
	4'b1111: F <= 2'b10;
	endcase
endmodule